-- FA_TB
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FA_TB IS
END FA_TB;

ARCHITECTURE HB OF FA_TB IS

	COMPONENT HB_FA
		PORT (
			A, B, CIN: IN BIT;
			S, COUT: OUT BIT
		);

	END COMPONENT;

	SIGNAL A: BIT := '0';
	SIGNAL B: BIT := '0';
	SIGNAL CIN: BIT := '0';
	SIGNAL S: BIT := '0';
	SIGNAL COUT: BIT := '0';

	BEGIN

		A <= '0', '0' AFTER 100NS, '1' AFTER 200NS, '1' AFTER 300NS, '1' AFTER 400NS;
		B <= '0', '0' AFTER 100NS, '0' AFTER 200NS, '1' AFTER 300NS, '1' AFTER 400NS;
		CIN <= '0', '1' AFTER 100NS, '0' AFTER 200NS, '0' AFTER 300NS, '1' AFTER 400NS;

	U1:HB_FA
	PORT MAP(
		A=>A,
		B=>B,
		CIN=>CIN,
		S=>S,
		COUT=>COUT
	);

END HB;