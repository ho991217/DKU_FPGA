-- TestBench of 8 to 3 encoder
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ENCODER_TB IS
END ENCODER_TB;


ARCHITECTURE HB OF ENCODER_TB IS

COMPONENT HB_ENCODER
PORT (
	I: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	O: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END COMPONENT;

SIGNAL I: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
SIGNAL O: STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";

BEGIN

I <= "00000001", "00000010" AFTER 100NS, "00000100" AFTER 200NS, "00001000" AFTER 300NS, "00010000" AFTER 400NS, "00100000" AFTER 500NS, "01000000" AFTER 600NS, "10000000" AFTER 700NS;

U1:HB_ENCODER
PORT MAP(
	I=>I,
	O=>O
);

END HB;
