-- TestBench of 3 to 8 decoder
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DECODER_TB IS
END DECODER_TB;

ARCHITECTURE HB OF DECODER_TB IS

COMPONENT HB_DECODER
PORT(
	A, B, C: IN STD_LOGIC;
	O: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;

SIGNAL A: STD_LOGIC := '0';
SIGNAL B: STD_LOGIC := '0';
SIGNAL C: STD_LOGIC := '0';
SIGNAL O: STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";

BEGIN

A <= '0', '1' AFTER 400NS;
B <= '0', '1' AFTER 200NS, '0' AFTER 400NS, '1' AFTER 600NS;
C <= '0', '1' AFTER 100NS, '0' AFTER 200NS, '1' AFTER 300NS, '0' AFTER 400NS, '1' AFTER 500NS, '0' AFTER 600NS, '0' AFTER 700NS, '1' AFTER 800NS;

U1:HB_DECODER
PORT MAP(
	A=>A,
	B=>B,
	C=>C,
	O=>O
);

END HB;