-- testbench
ENTITY EX_TB IS
END EX_TB;

ARCHITECTURE HB OF EX_TB IS

COMPONENT HB_EX
PORT(
	A, B: IN BIT;
	X: OUT BIT
);
END COMPONENT;

SIGNAL A: BIT := '0';
SIGNAL B: BIT := '0';
SIGNAL X: BIT := '0';

BEGIN

A <= '0', '1' AFTER 100NS, '0' AFTER 200NS, '1' AFTER 300NS; 
B <= '0', '0' AFTER 100NS, '1' AFTER 200NS, '1' AFTER 300NS;

U1:HB_EX
PORT MAP(
	A => A,
	B => B,
	X => X
);

END HB;